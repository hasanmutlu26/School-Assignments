magic
tech scmos
timestamp 1666631494
<< nwell >>
rect -17 18 43 28
<< polysilicon >>
rect -12 25 -10 27
rect -4 25 -2 27
rect 4 25 6 27
rect 20 25 22 27
rect 28 25 30 27
rect 36 25 38 27
rect -12 11 -10 21
rect -4 15 -2 21
rect 4 19 6 21
rect 20 19 22 21
rect 4 17 10 19
rect -4 13 6 15
rect -12 9 2 11
rect 0 6 2 9
rect 4 6 6 13
rect 8 6 10 17
rect 16 17 22 19
rect 16 6 18 17
rect 28 15 30 21
rect 20 13 30 15
rect 20 6 22 13
rect 36 11 38 21
rect 28 9 38 11
rect 28 6 30 9
rect 0 0 2 2
rect 4 0 6 2
rect 8 0 10 2
rect 16 0 18 2
rect 20 0 22 2
rect 28 0 30 2
<< ndiffusion >>
rect -1 2 0 6
rect 2 2 4 6
rect 6 2 8 6
rect 10 2 11 6
rect 15 2 16 6
rect 18 2 20 6
rect 22 2 23 6
rect 27 2 28 6
rect 30 2 31 6
<< pdiffusion >>
rect -13 21 -12 25
rect -10 21 -9 25
rect -5 21 -4 25
rect -2 21 -1 25
rect 3 21 4 25
rect 6 21 7 25
rect 19 21 20 25
rect 22 21 23 25
rect 27 21 28 25
rect 30 21 31 25
rect 35 21 36 25
rect 38 21 39 25
<< metal1 >>
rect -17 34 3 37
rect -17 25 -13 34
rect -1 25 3 34
rect 15 28 35 31
rect 15 25 19 28
rect 31 25 35 28
rect -9 18 -5 21
rect 7 18 11 21
rect 23 18 27 21
rect -9 15 27 18
rect 39 12 43 21
rect 11 9 43 12
rect 11 6 15 9
rect 31 6 35 9
rect -5 -1 -1 2
rect 23 -1 27 2
rect -5 -4 27 -1
<< ntransistor >>
rect 0 2 2 6
rect 4 2 6 6
rect 8 2 10 6
rect 16 2 18 6
rect 20 2 22 6
rect 28 2 30 6
<< ptransistor >>
rect -12 21 -10 25
rect -4 21 -2 25
rect 4 21 6 25
rect 20 21 22 25
rect 28 21 30 25
rect 36 21 38 25
<< ndcontact >>
rect -5 2 -1 6
rect 11 2 15 6
rect 23 2 27 6
rect 31 2 35 6
<< pdcontact >>
rect -17 21 -13 25
rect -9 21 -5 25
rect -1 21 3 25
rect 7 21 11 25
rect 15 21 19 25
rect 23 21 27 25
rect 31 21 35 25
rect 39 21 43 25
<< end >>
