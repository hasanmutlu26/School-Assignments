module _64bit_2x1MUX (result, A, B, control);
input [63:0] A, B;
input control;
output [63:0] result;

wire [63:0] and1, and2;

and (and1[0], A[0], ~control);
and (and1[1], A[1], ~control);
and (and1[2], A[2], ~control);
and (and1[3], A[3], ~control);
and (and1[4], A[4], ~control);
and (and1[5], A[5], ~control);
and (and1[6], A[6], ~control);
and (and1[7], A[7], ~control);
and (and1[8], A[8], ~control);
and (and1[9], A[9], ~control);
and (and1[10], A[10], ~control);
and (and1[11], A[11], ~control);
and (and1[12], A[12], ~control);
and (and1[13], A[13], ~control);
and (and1[14], A[14], ~control);
and (and1[15], A[15], ~control);
and (and1[16], A[16], ~control);
and (and1[17], A[17], ~control);
and (and1[18], A[18], ~control);
and (and1[19], A[19], ~control);
and (and1[20], A[20], ~control);
and (and1[21], A[21], ~control);
and (and1[22], A[22], ~control);
and (and1[23], A[23], ~control);
and (and1[24], A[24], ~control);
and (and1[25], A[25], ~control);
and (and1[26], A[26], ~control);
and (and1[27], A[27], ~control);
and (and1[28], A[28], ~control);
and (and1[29], A[29], ~control);
and (and1[30], A[30], ~control);
and (and1[31], A[31], ~control);
and (and1[32], A[32], ~control);
and (and1[33], A[33], ~control);
and (and1[34], A[34], ~control);
and (and1[35], A[35], ~control);
and (and1[36], A[36], ~control);
and (and1[37], A[37], ~control);
and (and1[38], A[38], ~control);
and (and1[39], A[39], ~control);
and (and1[40], A[40], ~control);
and (and1[41], A[41], ~control);
and (and1[42], A[42], ~control);
and (and1[43], A[43], ~control);
and (and1[44], A[44], ~control);
and (and1[45], A[45], ~control);
and (and1[46], A[46], ~control);
and (and1[47], A[47], ~control);
and (and1[48], A[48], ~control);
and (and1[49], A[49], ~control);
and (and1[50], A[50], ~control);
and (and1[51], A[51], ~control);
and (and1[52], A[52], ~control);
and (and1[53], A[53], ~control);
and (and1[54], A[54], ~control);
and (and1[55], A[55], ~control);
and (and1[56], A[56], ~control);
and (and1[57], A[57], ~control);
and (and1[58], A[58], ~control);
and (and1[59], A[59], ~control);
and (and1[60], A[60], ~control);
and (and1[61], A[61], ~control);
and (and1[62], A[62], ~control);
and (and1[63], A[63], ~control);

and (and2[0], B[0], control);
and (and2[1], B[1], control);
and (and2[2], B[2], control);
and (and2[3], B[3], control);
and (and2[4], B[4], control);
and (and2[5], B[5], control);
and (and2[6], B[6], control);
and (and2[7], B[7], control);
and (and2[8], B[8], control);
and (and2[9], B[9], control);
and (and2[10], B[10], control);
and (and2[11], B[11], control);
and (and2[12], B[12], control);
and (and2[13], B[13], control);
and (and2[14], B[14], control);
and (and2[15], B[15], control);
and (and2[16], B[16], control);
and (and2[17], B[17], control);
and (and2[18], B[18], control);
and (and2[19], B[19], control);
and (and2[20], B[20], control);
and (and2[21], B[21], control);
and (and2[22], B[22], control);
and (and2[23], B[23], control);
and (and2[24], B[24], control);
and (and2[25], B[25], control);
and (and2[26], B[26], control);
and (and2[27], B[27], control);
and (and2[28], B[28], control);
and (and2[29], B[29], control);
and (and2[30], B[30], control);
and (and2[31], B[31], control);
and (and2[32], B[32], control);
and (and2[33], B[33], control);
and (and2[34], B[34], control);
and (and2[35], B[35], control);
and (and2[36], B[36], control);
and (and2[37], B[37], control);
and (and2[38], B[38], control);
and (and2[39], B[39], control);
and (and2[40], B[40], control);
and (and2[41], B[41], control);
and (and2[42], B[42], control);
and (and2[43], B[43], control);
and (and2[44], B[44], control);
and (and2[45], B[45], control);
and (and2[46], B[46], control);
and (and2[47], B[47], control);
and (and2[48], B[48], control);
and (and2[49], B[49], control);
and (and2[50], B[50], control);
and (and2[51], B[51], control);
and (and2[52], B[52], control);
and (and2[53], B[53], control);
and (and2[54], B[54], control);
and (and2[55], B[55], control);
and (and2[56], B[56], control);
and (and2[57], B[57], control);
and (and2[58], B[58], control);
and (and2[59], B[59], control);
and (and2[60], B[60], control);
and (and2[61], B[61], control);
and (and2[62], B[62], control);
and (and2[63], B[63], control);

or (result[0], and1[0], and2[0]);
or (result[1], and1[1], and2[1]);
or (result[2], and1[2], and2[2]);
or (result[3], and1[3], and2[3]);
or (result[4], and1[4], and2[4]);
or (result[5], and1[5], and2[5]);
or (result[6], and1[6], and2[6]);
or (result[7], and1[7], and2[7]);
or (result[8], and1[8], and2[8]);
or (result[9], and1[9], and2[9]);
or (result[10], and1[10], and2[10]);
or (result[11], and1[11], and2[11]);
or (result[12], and1[12], and2[12]);
or (result[13], and1[13], and2[13]);
or (result[14], and1[14], and2[14]);
or (result[15], and1[15], and2[15]);
or (result[16], and1[16], and2[16]);
or (result[17], and1[17], and2[17]);
or (result[18], and1[18], and2[18]);
or (result[19], and1[19], and2[19]);
or (result[20], and1[20], and2[20]);
or (result[21], and1[21], and2[21]);
or (result[22], and1[22], and2[22]);
or (result[23], and1[23], and2[23]);
or (result[24], and1[24], and2[24]);
or (result[25], and1[25], and2[25]);
or (result[26], and1[26], and2[26]);
or (result[27], and1[27], and2[27]);
or (result[28], and1[28], and2[28]);
or (result[29], and1[29], and2[29]);
or (result[30], and1[30], and2[30]);
or (result[31], and1[31], and2[31]);
or (result[32], and1[32], and2[32]);
or (result[33], and1[33], and2[33]);
or (result[34], and1[34], and2[34]);
or (result[35], and1[35], and2[35]);
or (result[36], and1[36], and2[36]);
or (result[37], and1[37], and2[37]);
or (result[38], and1[38], and2[38]);
or (result[39], and1[39], and2[39]);
or (result[40], and1[40], and2[40]);
or (result[41], and1[41], and2[41]);
or (result[42], and1[42], and2[42]);
or (result[43], and1[43], and2[43]);
or (result[44], and1[44], and2[44]);
or (result[45], and1[45], and2[45]);
or (result[46], and1[46], and2[46]);
or (result[47], and1[47], and2[47]);
or (result[48], and1[48], and2[48]);
or (result[49], and1[49], and2[49]);
or (result[50], and1[50], and2[50]);
or (result[51], and1[51], and2[51]);
or (result[52], and1[52], and2[52]);
or (result[53], and1[53], and2[53]);
or (result[54], and1[54], and2[54]);
or (result[55], and1[55], and2[55]);
or (result[56], and1[56], and2[56]);
or (result[57], and1[57], and2[57]);
or (result[58], and1[58], and2[58]);
or (result[59], and1[59], and2[59]);
or (result[60], and1[60], and2[60]);
or (result[61], and1[61], and2[61]);
or (result[62], and1[62], and2[62]);
or (result[63], and1[63], and2[63]);

endmodule