magic
tech scmos
timestamp 1671278806
<< nwell >>
rect 128 98 135 118
<< metal1 >>
rect -1 116 0 120
rect 128 116 133 120
rect -1 57 0 61
rect 129 57 134 61
rect 262 57 263 61
rect -1 49 0 53
rect -1 32 4 36
rect -1 0 0 4
rect 129 0 134 4
<< m2contact >>
rect 4 31 9 36
<< metal2 >>
rect 136 36 140 51
rect 9 32 140 36
use xor2  xor2_1
timestamp 1671278367
transform 1 0 133 0 1 0
box -1 0 129 120
use xor2  xor2_0
timestamp 1671278367
transform 1 0 1 0 1 0
box -1 0 129 120
<< labels >>
rlabel metal1 0 32 0 36 3 C
rlabel metal1 0 57 0 61 3 A
rlabel metal1 0 49 0 53 3 B
rlabel metal1 0 0 0 4 2 gnd!
rlabel metal1 0 116 0 120 4 vdd!
rlabel metal1 262 57 262 61 7 Z
<< end >>
