module _32bit_8x1MUX_testbench();
reg [31:0] A,B,C,D,E,F,G,H;
reg [2:0] control;
wire [31:0] result;

_32bit_8x1MUX g0 (result, A,B,C,D,E,F,G,H,control);

initial begin
A = 32'b0000_0000_0000_0000_0000_0000_0000_1111;
B = 32'b0000_0000_0000_0000_0000_0000_1111_0000;
C = 32'b0000_0000_0000_0000_0000_1111_0000_0000;
D = 32'b0000_0000_0000_0000_1111_0000_0000_0000;
E = 32'b0000_0000_0000_1111_0000_0000_0000_0000;
F = 32'b0000_0000_1111_0000_0000_0000_0000_0000;
G = 32'b0000_1111_0000_0000_0000_0000_0000_0000;
H = 32'b1111_0000_0000_0000_0000_0000_0000_0000;

control = 3'b000;
#20;
control = 3'b001;
#20;
control = 3'b010;
#20;
control = 3'b011;
#20;
control = 3'b100;
#20;
control = 3'b101;
#20;
control = 3'b110;
#20;
control = 3'b111;
#20;

end

endmodule
