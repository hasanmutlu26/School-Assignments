magic
tech scmos
timestamp 1669032272
<< ntransistor >>
rect 5 6 7 10
rect 11 6 13 10
rect 19 6 21 10
rect 25 6 27 10
<< ptransistor >>
rect 5 30 7 34
rect 13 30 15 34
rect 29 30 31 34
rect 37 30 39 34
<< ndiffusion >>
rect 4 6 5 10
rect 7 6 11 10
rect 13 6 14 10
rect 18 6 19 10
rect 21 6 25 10
rect 27 6 28 10
<< pdiffusion >>
rect 4 30 5 34
rect 7 30 8 34
rect 12 30 13 34
rect 15 30 16 34
rect 28 30 29 34
rect 31 30 32 34
rect 36 30 37 34
rect 39 30 40 34
<< ndcontact >>
rect 0 6 4 10
rect 14 6 18 10
rect 28 6 32 10
<< pdcontact >>
rect 0 30 4 34
rect 8 30 12 34
rect 16 30 20 34
rect 24 30 28 34
rect 32 30 36 34
rect 40 30 44 34
<< polysilicon >>
rect 5 34 7 37
rect 13 34 15 37
rect 29 34 31 37
rect 37 34 39 37
rect 5 10 7 30
rect 13 29 15 30
rect 29 29 31 30
rect 11 27 15 29
rect 19 27 31 29
rect 11 10 13 27
rect 19 10 21 27
rect 37 22 39 30
rect 25 20 39 22
rect 25 10 27 20
rect 5 3 7 6
rect 11 3 13 6
rect 19 3 21 6
rect 25 3 27 6
<< metal1 >>
rect 0 38 20 41
rect 0 34 4 38
rect 16 34 20 38
rect 24 38 44 41
rect 24 34 28 38
rect 40 34 44 38
rect 8 26 12 30
rect 32 26 36 30
rect 8 22 36 26
rect 40 18 44 30
rect 14 14 44 18
rect 14 10 18 14
rect 0 2 4 6
rect 28 2 32 6
rect 0 -2 32 2
<< labels >>
rlabel metal1 0 -2 0 2 2 gnd!
rlabel space 0 38 0 42 4 vdd!
rlabel metal1 44 14 44 18 7 Y
rlabel polysilicon 5 3 7 3 1 A
rlabel polysilicon 11 3 13 3 1 B
rlabel polysilicon 19 3 21 3 1 C
rlabel polysilicon 25 3 27 3 1 D
<< end >>
