module _64bit_shiftRight(result, A, control);
input [63:0] A;
input control;
output [63:0] result;


_1bit_2x1MUX g1 (result[0], A[0], A[1], control);
_1bit_2x1MUX g2 (result[1], A[1], A[2], control);
_1bit_2x1MUX g3 (result[2], A[2], A[3], control);
_1bit_2x1MUX g4 (result[3], A[3], A[4], control);
_1bit_2x1MUX g5 (result[4], A[4], A[5], control);
_1bit_2x1MUX g6 (result[5], A[5], A[6], control);
_1bit_2x1MUX g7 (result[6], A[6], A[7], control);
_1bit_2x1MUX g8 (result[7], A[7], A[8], control);
_1bit_2x1MUX g9 (result[8], A[8], A[9], control);
_1bit_2x1MUX g10 (result[9], A[9], A[10], control);
_1bit_2x1MUX g11 (result[10], A[10], A[11], control);
_1bit_2x1MUX g12 (result[11], A[11], A[12], control);
_1bit_2x1MUX g13 (result[12], A[12], A[13], control);
_1bit_2x1MUX g14 (result[13], A[13], A[14], control);
_1bit_2x1MUX g15 (result[14], A[14], A[15], control);
_1bit_2x1MUX g16 (result[15], A[15], A[16], control);
_1bit_2x1MUX g17 (result[16], A[16], A[17], control);
_1bit_2x1MUX g18 (result[17], A[17], A[18], control);
_1bit_2x1MUX g19 (result[18], A[18], A[19], control);
_1bit_2x1MUX g20 (result[19], A[19], A[20], control);
_1bit_2x1MUX g21 (result[20], A[20], A[21], control);
_1bit_2x1MUX g22 (result[21], A[21], A[22], control);
_1bit_2x1MUX g23 (result[22], A[22], A[23], control);
_1bit_2x1MUX g24 (result[23], A[23], A[24], control);
_1bit_2x1MUX g25 (result[24], A[24], A[25], control);
_1bit_2x1MUX g26 (result[25], A[25], A[26], control);
_1bit_2x1MUX g27 (result[26], A[26], A[27], control);
_1bit_2x1MUX g28 (result[27], A[27], A[28], control);
_1bit_2x1MUX g29 (result[28], A[28], A[29], control);
_1bit_2x1MUX g30 (result[29], A[29], A[30], control);
_1bit_2x1MUX g31 (result[30], A[30], A[31], control);
_1bit_2x1MUX g32 (result[31], A[31], A[32], control);
_1bit_2x1MUX g33 (result[32], A[32], A[33], control);
_1bit_2x1MUX g34 (result[33], A[33], A[34], control);
_1bit_2x1MUX g35 (result[34], A[34], A[35], control);
_1bit_2x1MUX g36 (result[35], A[35], A[36], control);
_1bit_2x1MUX g37 (result[36], A[36], A[37], control);
_1bit_2x1MUX g38 (result[37], A[37], A[38], control);
_1bit_2x1MUX g39 (result[38], A[38], A[39], control);
_1bit_2x1MUX g40 (result[39], A[39], A[40], control);
_1bit_2x1MUX g41 (result[40], A[40], A[41], control);
_1bit_2x1MUX g42 (result[41], A[41], A[42], control);
_1bit_2x1MUX g43 (result[42], A[42], A[43], control);
_1bit_2x1MUX g44 (result[43], A[43], A[44], control);
_1bit_2x1MUX g45 (result[44], A[44], A[45], control);
_1bit_2x1MUX g46 (result[45], A[45], A[46], control);
_1bit_2x1MUX g47 (result[46], A[46], A[47], control);
_1bit_2x1MUX g48 (result[47], A[47], A[48], control);
_1bit_2x1MUX g49 (result[48], A[48], A[49], control);
_1bit_2x1MUX g50 (result[49], A[49], A[50], control);
_1bit_2x1MUX g51 (result[50], A[50], A[51], control);
_1bit_2x1MUX g52 (result[51], A[51], A[52], control);
_1bit_2x1MUX g53 (result[52], A[52], A[53], control);
_1bit_2x1MUX g54 (result[53], A[53], A[54], control);
_1bit_2x1MUX g55 (result[54], A[54], A[55], control);
_1bit_2x1MUX g56 (result[55], A[55], A[56], control);
_1bit_2x1MUX g57 (result[56], A[56], A[57], control);
_1bit_2x1MUX g58 (result[57], A[57], A[58], control);
_1bit_2x1MUX g59 (result[58], A[58], A[59], control);
_1bit_2x1MUX g60 (result[59], A[59], A[60], control);
_1bit_2x1MUX g61 (result[60], A[60], A[61], control);
_1bit_2x1MUX g62 (result[61], A[61], A[62], control);
_1bit_2x1MUX g63 (result[62], A[62], A[63], control);
_1bit_2x1MUX g64 (result[63], A[63], 1'b0, control);

endmodule