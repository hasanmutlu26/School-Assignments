magic
tech scmos
timestamp 1669031839
<< ntransistor >>
rect 5 8 7 12
<< ptransistor >>
rect 5 31 7 35
<< ndiffusion >>
rect 4 8 5 12
rect 7 8 8 12
<< pdiffusion >>
rect 4 31 5 35
rect 7 31 8 35
<< ndcontact >>
rect 0 8 4 12
rect 8 8 12 12
<< pdcontact >>
rect 0 31 4 35
rect 8 31 12 35
<< polysilicon >>
rect 5 35 7 38
rect 5 12 7 31
rect 5 5 7 8
<< metal1 >>
rect 0 39 12 43
rect 0 35 4 39
rect 8 12 12 31
rect 0 4 4 8
rect 0 0 12 4
<< labels >>
rlabel metal1 12 19 12 23 7 Y
rlabel polysilicon 5 5 7 5 1 A
rlabel metal1 0 39 0 43 4 vdd!
rlabel metal1 0 0 0 4 2 gnd!
<< end >>
