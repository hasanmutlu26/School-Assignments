module _64bit_register (value, data, clk);
input [63:0] data;
input clk;
output [63:0] value;

DFlipFlop g0 (value[0], ,data[0], clk);
DFlipFlop g1 (value[1], ,data[1], clk);
DFlipFlop g2 (value[2], ,data[2], clk);
DFlipFlop g3 (value[3], ,data[3], clk);
DFlipFlop g4 (value[4], ,data[4], clk);
DFlipFlop g5 (value[5], ,data[5], clk);
DFlipFlop g6 (value[6], ,data[6], clk);
DFlipFlop g7 (value[7], ,data[7], clk);
DFlipFlop g8 (value[8], ,data[8], clk);
DFlipFlop g9 (value[9], ,data[9], clk);
DFlipFlop g10 (value[10], ,data[10], clk);
DFlipFlop g11 (value[11], ,data[11], clk);
DFlipFlop g12 (value[12], ,data[12], clk);
DFlipFlop g13 (value[13], ,data[13], clk);
DFlipFlop g14 (value[14], ,data[14], clk);
DFlipFlop g15 (value[15], ,data[15], clk);
DFlipFlop g16 (value[16], ,data[16], clk);
DFlipFlop g17 (value[17], ,data[17], clk);
DFlipFlop g18 (value[18], ,data[18], clk);
DFlipFlop g19 (value[19], ,data[19], clk);
DFlipFlop g20 (value[20], ,data[20], clk);
DFlipFlop g21 (value[21], ,data[21], clk);
DFlipFlop g22 (value[22], ,data[22], clk);
DFlipFlop g23 (value[23], ,data[23], clk);
DFlipFlop g24 (value[24], ,data[24], clk);
DFlipFlop g25 (value[25], ,data[25], clk);
DFlipFlop g26 (value[26], ,data[26], clk);
DFlipFlop g27 (value[27], ,data[27], clk);
DFlipFlop g28 (value[28], ,data[28], clk);
DFlipFlop g29 (value[29], ,data[29], clk);
DFlipFlop g30 (value[30], ,data[30], clk);
DFlipFlop g31 (value[31], ,data[31], clk);
DFlipFlop g32 (value[32], ,data[32], clk);
DFlipFlop g33 (value[33], ,data[33], clk);
DFlipFlop g34 (value[34], ,data[34], clk);
DFlipFlop g35 (value[35], ,data[35], clk);
DFlipFlop g36 (value[36], ,data[36], clk);
DFlipFlop g37 (value[37], ,data[37], clk);
DFlipFlop g38 (value[38], ,data[38], clk);
DFlipFlop g39 (value[39], ,data[39], clk);
DFlipFlop g40 (value[40], ,data[40], clk);
DFlipFlop g41 (value[41], ,data[41], clk);
DFlipFlop g42 (value[42], ,data[42], clk);
DFlipFlop g43 (value[43], ,data[43], clk);
DFlipFlop g44 (value[44], ,data[44], clk);
DFlipFlop g45 (value[45], ,data[45], clk);
DFlipFlop g46 (value[46], ,data[46], clk);
DFlipFlop g47 (value[47], ,data[47], clk);
DFlipFlop g48 (value[48], ,data[48], clk);
DFlipFlop g49 (value[49], ,data[49], clk);
DFlipFlop g50 (value[50], ,data[50], clk);
DFlipFlop g51 (value[51], ,data[51], clk);
DFlipFlop g52 (value[52], ,data[52], clk);
DFlipFlop g53 (value[53], ,data[53], clk);
DFlipFlop g54 (value[54], ,data[54], clk);
DFlipFlop g55 (value[55], ,data[55], clk);
DFlipFlop g56 (value[56], ,data[56], clk);
DFlipFlop g57 (value[57], ,data[57], clk);
DFlipFlop g58 (value[58], ,data[58], clk);
DFlipFlop g59 (value[59], ,data[59], clk);
DFlipFlop g60 (value[60], ,data[60], clk);
DFlipFlop g61 (value[61], ,data[61], clk);
DFlipFlop g62 (value[62], ,data[62], clk);
DFlipFlop g63 (value[63], ,data[63], clk);

endmodule