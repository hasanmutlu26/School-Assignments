library verilog;
use verilog.vl_types.all;
entity \_32bit_SLT_testbench\ is
end \_32bit_SLT_testbench\;
